<svg xmlns="http://www.w3.org/2000/svg" width="480" height="330" class="">
    <defs>
        <style/>
    </defs>
    <style>@keyframes animation-gauge{0%{stroke-dasharray:0 329}}@keyframes animation-rainbow{0%,to{color:#7f00ff;fill:#7f00ff}14%{color:#a933ff;fill:#a933ff}29%{color:#007fff;fill:#007fff}43%{color:#00ff7f;fill:#00ff7f}57%{color:#ff0;fill:#ff0}71%{color:#ff7f00;fill:#ff7f00}86%{color:red;fill:red}}svg{font-family:-apple-system,BlinkMacSystemFont,Segoe UI,Helvetica,Arial,sans-serif,Apple Color Emoji,Segoe UI Emoji;color:#777}h2,h3{margin:8px 0 2px;padding:0;color:#0366d6;font-weight:400}h2 svg,h3 svg{fill:currentColor}h2{font-size:16px}h3,svg{font-size:14px}section&gt;.field{margin-left:5px;margin-right:5px}.field{display:flex;align-items:center;margin-bottom:2px;white-space:nowrap}.field svg{margin:0 8px;fill:#959da5;flex-shrink:0}.row{display:flex;flex-wrap:wrap}.row section{flex:1 1 0}.calendar.field{margin:4px 0 4px 7px}.calendar .day{outline:1px solid rgba(27,31,35,.04);outline-offset:-1px}svg.calendar{margin-left:13px;margin-top:4px}:root{--color-calendar-graph-day-bg:#ebedf0;--color-calendar-graph-day-border:rgba(27,31,35,0.06);--color-calendar-graph-day-L1-bg:#9be9a8;--color-calendar-graph-day-L2-bg:#40c463;--color-calendar-graph-day-L3-bg:#30a14e;--color-calendar-graph-day-L4-bg:#216e39;--color-calendar-halloween-graph-day-L1-bg:#ffee4a;--color-calendar-halloween-graph-day-L2-bg:#ffc501;--color-calendar-halloween-graph-day-L3-bg:#fe9600;--color-calendar-halloween-graph-day-L4-bg:#03001c;--color-calendar-winter-graph-day-L1-bg:#0a3069;--color-calendar-winter-graph-day-L2-bg:#0969da;--color-calendar-winter-graph-day-L3-bg:#54aeff;--color-calendar-winter-graph-day-L4-bg:#b6e3ff;--color-calendar-graph-day-L4-border:rgba(27,31,35,0.06);--color-calendar-graph-day-L3-border:rgba(27,31,35,0.06);--color-calendar-graph-day-L2-border:rgba(27,31,35,0.06);--color-calendar-graph-day-L1-border:rgba(27,31,35,0.06)}#metrics-end{width:100%}</style>
    <style/>
    <foreignObject x="0" y="0" width="100%" height="100%">
        <div xmlns="http://www.w3.org/1999/xhtml" xmlns:xlink="http://www.w3.org/1999/xlink" class="items-wrapper">
            <section>
                <h2 class="field">
                    <svg xmlns="http://www.w3.org/2000/svg" viewBox="0 0 16 16" width="16" height="16">
                        <path fill-rule="evenodd" d="M4.75 0a.75.75 0 01.75.75V2h5V.75a.75.75 0 011.5 0V2h1.25c.966 0 1.75.784 1.75 1.75v10.5A1.75 1.75 0 0113.25 16H2.75A1.75 1.75 0 011 14.25V3.75C1 2.784 1.784 2 2.75 2H4V.75A.75.75 0 014.75 0zm0 3.5h8.5a.25.25 0 01.25.25V6h-11V3.75a.25.25 0 01.25-.25h2zm-2.25 4v6.75c0 .138.112.25.25.25h10.5a.25.25 0 00.25-.25V7.5h-11z"/>
                    </svg>
                    Contributions calendar
                </h2>
                <div class="row">
                    <section>
                    </section>
                    <section>
                        <h3 class="field">
                            <svg xmlns="http://www.w3.org/2000/svg" viewBox="0 0 16 16" width="16" height="16">
                                <path fill-rule="evenodd" d="M7.75 14A1.75 1.75 0 016 12.25v-8.5C6 2.784 6.784 2 7.75 2h6.5c.966 0 1.75.784 1.75 1.75v8.5A1.75 1.75 0 0114.25 14h-6.5zm-.25-1.75c0 .138.112.25.25.25h6.5a.25.25 0 00.25-.25v-8.5a.25.25 0 00-.25-.25h-6.5a.25.25 0 00-.25.25v8.5zM4.9 3.508a.75.75 0 01-.274 1.025.25.25 0 00-.126.217v6.5a.25.25 0 00.126.217.75.75 0 01-.752 1.298A1.75 1.75 0 013 11.25v-6.5c0-.649.353-1.214.874-1.516a.75.75 0 011.025.274zM1.625 5.533a.75.75 0 10-.752-1.299A1.75 1.75 0 000 5.75v4.5c0 .649.353 1.214.874 1.515a.75.75 0 10.752-1.298.25.25 0 01-.126-.217v-4.5a.25.25 0 01.126-.217z"/>
                            </svg>
                            Commits streaks
                        </h3>
                        <div class="field">
                            <svg xmlns="http://www.w3.org/2000/svg" viewBox="0 0 16 16" width="16" height="16">
                                <path fill-rule="evenodd" d="M7.998 14.5c2.832 0 5-1.98 5-4.5 0-1.463-.68-2.19-1.879-3.383l-.036-.037c-1.013-1.008-2.3-2.29-2.834-4.434-.322.256-.63.579-.864.953-.432.696-.621 1.58-.046 2.73.473.947.67 2.284-.278 3.232-.61.61-1.545.84-2.403.633a2.788 2.788 0 01-1.436-.874A3.21 3.21 0 003 10c0 2.53 2.164 4.5 4.998 4.5zM9.533.753C9.496.34 9.16.009 8.77.146 7.035.75 4.34 3.187 5.997 6.5c.344.689.285 1.218.003 1.5-.419.419-1.54.487-2.04-.832-.173-.454-.659-.762-1.035-.454C2.036 7.44 1.5 8.702 1.5 10c0 3.512 2.998 6 6.498 6s6.5-2.5 6.5-6c0-2.137-1.128-3.26-2.312-4.438-1.19-1.184-2.436-2.425-2.653-4.81z"/>
                            </svg>
                            Current streak 6 days
                        </div>
                        <div class="field">
                            <svg xmlns="http://www.w3.org/2000/svg" viewBox="0 0 16 16" width="16" height="16">
                                <path d="M8.5.75a.75.75 0 00-1.5 0v5.19L4.391 3.33a.75.75 0 10-1.06 1.061L5.939 7H.75a.75.75 0 000 1.5h5.19l-2.61 2.609a.75.75 0 101.061 1.06L7 9.561v5.189a.75.75 0 001.5 0V9.56l2.609 2.61a.75.75 0 101.06-1.061L9.561 8.5h5.189a.75.75 0 000-1.5H9.56l2.61-2.609a.75.75 0 00-1.061-1.06L8.5 5.939V.75z"/>
                            </svg>
                            Best streak 35 days
                        </div>
                        <h3 class="field">
                            <svg xmlns="http://www.w3.org/2000/svg" viewBox="0 0 16 16" width="16" height="16">
                                <path fill-rule="evenodd" d="M10.5 7.75a2.5 2.5 0 11-5 0 2.5 2.5 0 015 0zm1.43.75a4.002 4.002 0 01-7.86 0H.75a.75.75 0 110-1.5h3.32a4.001 4.001 0 017.86 0h3.32a.75.75 0 110 1.5h-3.32z"/>
                            </svg>
                            Commits per day
                        </h3>
                        <div class="field">
                            <svg xmlns="http://www.w3.org/2000/svg" viewBox="0 0 16 16" width="16" height="16">
                                <path d="M7.823 1.677L4.927 4.573A.25.25 0 005.104 5H7.25v3.236a.75.75 0 101.5 0V5h2.146a.25.25 0 00.177-.427L8.177 1.677a.25.25 0 00-.354 0zM13.75 11a.75.75 0 000 1.5h.5a.75.75 0 000-1.5h-.5zm-3.75.75a.75.75 0 01.75-.75h.5a.75.75 0 010 1.5h-.5a.75.75 0 01-.75-.75zM7.75 11a.75.75 0 000 1.5h.5a.75.75 0 000-1.5h-.5zM4 11.75a.75.75 0 01.75-.75h.5a.75.75 0 010 1.5h-.5a.75.75 0 01-.75-.75zM1.75 11a.75.75 0 000 1.5h.5a.75.75 0 000-1.5h-.5z"/>
                            </svg>
                            Highest in a day at 57
                        </div>
                        <div class="field">
                            <svg xmlns="http://www.w3.org/2000/svg" viewBox="0 0 16 16" width="16" height="16">
                                <path d="M10.896 2H8.75V.75a.75.75 0 00-1.5 0V2H5.104a.25.25 0 00-.177.427l2.896 2.896a.25.25 0 00.354 0l2.896-2.896A.25.25 0 0010.896 2zM8.75 15.25a.75.75 0 01-1.5 0V14H5.104a.25.25 0 01-.177-.427l2.896-2.896a.25.25 0 01.354 0l2.896 2.896a.25.25 0 01-.177.427H8.75v1.25zm-6.5-6.5a.75.75 0 000-1.5h-.5a.75.75 0 000 1.5h.5zM6 8a.75.75 0 01-.75.75h-.5a.75.75 0 010-1.5h.5A.75.75 0 016 8zm2.25.75a.75.75 0 000-1.5h-.5a.75.75 0 000 1.5h.5zM12 8a.75.75 0 01-.75.75h-.5a.75.75 0 010-1.5h.5A.75.75 0 0112 8zm2.25.75a.75.75 0 000-1.5h-.5a.75.75 0 000 1.5h.5z"/>
                            </svg>
                            Average per day at ~6.15
                        </div>
                    </section>
                </div>
                <svg version="1.1" xmlns="http://www.w3.org/2000/svg" style="margin-top: -130px;" viewBox="0,0 480,270">
                    <filter id="brightness1">
                        <feComponentTransfer>
                            <feFuncR type="linear" slope="0.6"/>
                            <feFuncG type="linear" slope="0.6"/>
                            <feFuncB type="linear" slope="0.6"/>
                        </feComponentTransfer>
                    </filter>
                    <filter id="brightness2">
                        <feComponentTransfer>
                            <feFuncR type="linear" slope="0.19999999999999996"/>
                            <feFuncG type="linear" slope="0.19999999999999996"/>
                            <feFuncB type="linear" slope="0.19999999999999996"/>
                        </feComponentTransfer>
                    </filter>
                    <g transform="scale(4) translate(12, 0)">
                        <g transform="translate(0, 0)">
                            <g transform="translate(0, 5.578947368421053)">
                                <path fill="#40c463" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#40c463" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.4210526315789473 0,1.4210526315789473 z"/>
                                <path fill="#40c463" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.4210526315789473 1.7,2.4210526315789473 z"/>
                            </g>
                            <g transform="translate(-1.7, 6.684210526315789)">
                                <path fill="#9be9a8" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#9be9a8" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.3157894736842106 0,1.3157894736842106 z"/>
                                <path fill="#9be9a8" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.3157894736842106 1.7,2.3157894736842106 z"/>
                            </g>
                            <g transform="translate(-3.4, 6.842105263157896)">
                                <path fill="#216e39" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#216e39" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,3.1578947368421053 0,2.1578947368421053 z"/>
                                <path fill="#216e39" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,2.1578947368421053 1.7,3.1578947368421053 z"/>
                            </g>
                            <g transform="translate(-5.1, 8.157894736842106)">
                                <path fill="#30a14e" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#30a14e" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.8421052631578947 0,1.8421052631578947 z"/>
                                <path fill="#30a14e" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.8421052631578947 1.7,2.8421052631578947 z"/>
                            </g>
                            <g transform="translate(-6.8, 10)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-8.5, 11)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-10.2, 12)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                        </g>
                        <g transform="translate(1.7, 1)">
                            <g transform="translate(0, 6)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-1.7, 5.631578947368421)">
                                <path fill="#216e39" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#216e39" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,3.3684210526315788 0,2.3684210526315788 z"/>
                                <path fill="#216e39" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,2.3684210526315788 1.7,3.3684210526315788 z"/>
                            </g>
                            <g transform="translate(-3.4, 7.578947368421053)">
                                <path fill="#40c463" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#40c463" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.4210526315789473 0,1.4210526315789473 z"/>
                                <path fill="#40c463" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.4210526315789473 1.7,2.4210526315789473 z"/>
                            </g>
                            <g transform="translate(-5.1, 8.473684210526315)">
                                <path fill="#40c463" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#40c463" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.526315789473684 0,1.526315789473684 z"/>
                                <path fill="#40c463" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.526315789473684 1.7,2.526315789473684 z"/>
                            </g>
                            <g transform="translate(-6.8, 8.947368421052632)">
                                <path fill="#216e39" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#216e39" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,3.052631578947368 0,2.052631578947368 z"/>
                                <path fill="#216e39" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,2.052631578947368 1.7,3.052631578947368 z"/>
                            </g>
                            <g transform="translate(-8.5, 10.157894736842106)">
                                <path fill="#30a14e" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#30a14e" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.8421052631578947 0,1.8421052631578947 z"/>
                                <path fill="#30a14e" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.8421052631578947 1.7,2.8421052631578947 z"/>
                            </g>
                            <g transform="translate(-10.2, 12)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                        </g>
                        <g transform="translate(3.4, 2)">
                            <g transform="translate(0, 5.894736842105263)">
                                <path fill="#9be9a8" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#9be9a8" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.1052631578947367 0,1.1052631578947367 z"/>
                                <path fill="#9be9a8" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.1052631578947367 1.7,2.1052631578947367 z"/>
                            </g>
                            <g transform="translate(-1.7, 5.947368421052632)">
                                <path fill="#216e39" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#216e39" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,3.052631578947368 0,2.052631578947368 z"/>
                                <path fill="#216e39" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,2.052631578947368 1.7,3.052631578947368 z"/>
                            </g>
                            <g transform="translate(-3.4, 7.368421052631579)">
                                <path fill="#40c463" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#40c463" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.6315789473684212 0,1.631578947368421 z"/>
                                <path fill="#40c463" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.631578947368421 1.7,2.6315789473684212 z"/>
                            </g>
                            <g transform="translate(-5.1, 8.263157894736842)">
                                <path fill="#30a14e" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#30a14e" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.736842105263158 0,1.736842105263158 z"/>
                                <path fill="#30a14e" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.736842105263158 1.7,2.736842105263158 z"/>
                            </g>
                            <g transform="translate(-6.8, 9.578947368421053)">
                                <path fill="#40c463" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#40c463" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.4210526315789473 0,1.4210526315789473 z"/>
                                <path fill="#40c463" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.4210526315789473 1.7,2.4210526315789473 z"/>
                            </g>
                            <g transform="translate(-8.5, 10.473684210526315)">
                                <path fill="#40c463" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#40c463" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.526315789473684 0,1.526315789473684 z"/>
                                <path fill="#40c463" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.526315789473684 1.7,2.526315789473684 z"/>
                            </g>
                            <g transform="translate(-10.2, 12)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                        </g>
                        <g transform="translate(5.1, 3)">
                            <g transform="translate(0, 5.684210526315789)">
                                <path fill="#9be9a8" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#9be9a8" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.3157894736842106 0,1.3157894736842106 z"/>
                                <path fill="#9be9a8" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.3157894736842106 1.7,2.3157894736842106 z"/>
                            </g>
                            <g transform="translate(-1.7, 6.578947368421053)">
                                <path fill="#40c463" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#40c463" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.4210526315789473 0,1.4210526315789473 z"/>
                                <path fill="#40c463" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.4210526315789473 1.7,2.4210526315789473 z"/>
                            </g>
                            <g transform="translate(-3.4, 7.052631578947368)">
                                <path fill="#30a14e" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#30a14e" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.9473684210526314 0,1.9473684210526314 z"/>
                                <path fill="#30a14e" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.9473684210526314 1.7,2.9473684210526314 z"/>
                            </g>
                            <g transform="translate(-5.1, 7.947368421052632)">
                                <path fill="#216e39" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#216e39" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,3.052631578947368 0,2.052631578947368 z"/>
                                <path fill="#216e39" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,2.052631578947368 1.7,3.052631578947368 z"/>
                            </g>
                            <g transform="translate(-6.8, 9.68421052631579)">
                                <path fill="#9be9a8" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#9be9a8" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.3157894736842106 0,1.3157894736842106 z"/>
                                <path fill="#9be9a8" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.3157894736842106 1.7,2.3157894736842106 z"/>
                            </g>
                            <g transform="translate(-8.5, 9.631578947368421)">
                                <path fill="#216e39" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#216e39" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,3.3684210526315788 0,2.3684210526315788 z"/>
                                <path fill="#216e39" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,2.3684210526315788 1.7,3.3684210526315788 z"/>
                            </g>
                            <g transform="translate(-10.2, 11.368421052631579)">
                                <path fill="#40c463" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#40c463" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.6315789473684212 0,1.631578947368421 z"/>
                                <path fill="#40c463" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.631578947368421 1.7,2.6315789473684212 z"/>
                            </g>
                        </g>
                        <g transform="translate(6.8, 4)">
                            <g transform="translate(0, 6)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-1.7, 6.052631578947368)">
                                <path fill="#30a14e" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#30a14e" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.9473684210526314 0,1.9473684210526314 z"/>
                                <path fill="#30a14e" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.9473684210526314 1.7,2.9473684210526314 z"/>
                            </g>
                            <g transform="translate(-3.4, 6.7368421052631575)">
                                <path fill="#216e39" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#216e39" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,3.263157894736842 0,2.263157894736842 z"/>
                                <path fill="#216e39" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,2.263157894736842 1.7,3.263157894736842 z"/>
                            </g>
                            <g transform="translate(-5.1, 8.368421052631579)">
                                <path fill="#40c463" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#40c463" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.6315789473684212 0,1.631578947368421 z"/>
                                <path fill="#40c463" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.631578947368421 1.7,2.6315789473684212 z"/>
                            </g>
                            <g transform="translate(-6.8, 9.368421052631579)">
                                <path fill="#40c463" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#40c463" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.6315789473684212 0,1.631578947368421 z"/>
                                <path fill="#40c463" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.631578947368421 1.7,2.6315789473684212 z"/>
                            </g>
                            <g transform="translate(-8.5, 9.631578947368421)">
                                <path fill="#216e39" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#216e39" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,3.3684210526315788 0,2.3684210526315788 z"/>
                                <path fill="#216e39" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,2.3684210526315788 1.7,3.3684210526315788 z"/>
                            </g>
                            <g transform="translate(-10.2, 11.894736842105264)">
                                <path fill="#9be9a8" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#9be9a8" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.1052631578947367 0,1.1052631578947367 z"/>
                                <path fill="#9be9a8" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.1052631578947367 1.7,2.1052631578947367 z"/>
                            </g>
                        </g>
                        <g transform="translate(8.5, 5)">
                            <g transform="translate(0, 5.684210526315789)">
                                <path fill="#9be9a8" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#9be9a8" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.3157894736842106 0,1.3157894736842106 z"/>
                                <path fill="#9be9a8" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.3157894736842106 1.7,2.3157894736842106 z"/>
                            </g>
                            <g transform="translate(-1.7, 5.526315789473684)">
                                <path fill="#216e39" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#216e39" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,3.473684210526316 0,2.473684210526316 z"/>
                                <path fill="#216e39" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,2.473684210526316 1.7,3.473684210526316 z"/>
                            </g>
                            <g transform="translate(-3.4, 6.631578947368421)">
                                <path fill="#216e39" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#216e39" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,3.3684210526315788 0,2.3684210526315788 z"/>
                                <path fill="#216e39" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,2.3684210526315788 1.7,3.3684210526315788 z"/>
                            </g>
                            <g transform="translate(-5.1, 8.473684210526315)">
                                <path fill="#40c463" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#40c463" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.526315789473684 0,1.526315789473684 z"/>
                                <path fill="#40c463" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.526315789473684 1.7,2.526315789473684 z"/>
                            </g>
                            <g transform="translate(-6.8, 9.578947368421053)">
                                <path fill="#40c463" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#40c463" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.4210526315789473 0,1.4210526315789473 z"/>
                                <path fill="#40c463" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.4210526315789473 1.7,2.4210526315789473 z"/>
                            </g>
                            <g transform="translate(-8.5, 9.736842105263158)">
                                <path fill="#216e39" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#216e39" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,3.263157894736842 0,2.263157894736842 z"/>
                                <path fill="#216e39" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,2.263157894736842 1.7,3.263157894736842 z"/>
                            </g>
                            <g transform="translate(-10.2, 11.68421052631579)">
                                <path fill="#9be9a8" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#9be9a8" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.3157894736842106 0,1.3157894736842106 z"/>
                                <path fill="#9be9a8" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.3157894736842106 1.7,2.3157894736842106 z"/>
                            </g>
                        </g>
                        <g transform="translate(10.2, 6)">
                            <g transform="translate(0, 5.684210526315789)">
                                <path fill="#9be9a8" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#9be9a8" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.3157894736842106 0,1.3157894736842106 z"/>
                                <path fill="#9be9a8" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.3157894736842106 1.7,2.3157894736842106 z"/>
                            </g>
                            <g transform="translate(-1.7, 5.526315789473684)">
                                <path fill="#216e39" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#216e39" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,3.473684210526316 0,2.473684210526316 z"/>
                                <path fill="#216e39" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,2.473684210526316 1.7,3.473684210526316 z"/>
                            </g>
                            <g transform="translate(-3.4, 7.684210526315789)">
                                <path fill="#9be9a8" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#9be9a8" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.3157894736842106 0,1.3157894736842106 z"/>
                                <path fill="#9be9a8" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.3157894736842106 1.7,2.3157894736842106 z"/>
                            </g>
                            <g transform="translate(-5.1, 8.157894736842106)">
                                <path fill="#30a14e" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#30a14e" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.8421052631578947 0,1.8421052631578947 z"/>
                                <path fill="#30a14e" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.8421052631578947 1.7,2.8421052631578947 z"/>
                            </g>
                            <g transform="translate(-6.8, 9.263157894736842)">
                                <path fill="#40c463" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#40c463" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.736842105263158 0,1.736842105263158 z"/>
                                <path fill="#40c463" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.736842105263158 1.7,2.736842105263158 z"/>
                            </g>
                            <g transform="translate(-8.5, 10.263157894736842)">
                                <path fill="#40c463" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#40c463" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.736842105263158 0,1.736842105263158 z"/>
                                <path fill="#40c463" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.736842105263158 1.7,2.736842105263158 z"/>
                            </g>
                            <g transform="translate(-10.2, 11.789473684210527)">
                                <path fill="#9be9a8" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#9be9a8" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.2105263157894735 0,1.2105263157894737 z"/>
                                <path fill="#9be9a8" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.2105263157894737 1.7,2.2105263157894735 z"/>
                            </g>
                        </g>
                        <g transform="translate(11.9, 7)">
                            <g transform="translate(0, 6)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-1.7, 6.473684210526315)">
                                <path fill="#40c463" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#40c463" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.526315789473684 0,1.526315789473684 z"/>
                                <path fill="#40c463" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.526315789473684 1.7,2.526315789473684 z"/>
                            </g>
                            <g transform="translate(-3.4, 7.894736842105263)">
                                <path fill="#9be9a8" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#9be9a8" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.1052631578947367 0,1.1052631578947367 z"/>
                                <path fill="#9be9a8" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.1052631578947367 1.7,2.1052631578947367 z"/>
                            </g>
                            <g transform="translate(-5.1, 8.68421052631579)">
                                <path fill="#9be9a8" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#9be9a8" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.3157894736842106 0,1.3157894736842106 z"/>
                                <path fill="#9be9a8" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.3157894736842106 1.7,2.3157894736842106 z"/>
                            </g>
                            <g transform="translate(-6.8, 9.894736842105264)">
                                <path fill="#9be9a8" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#9be9a8" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.1052631578947367 0,1.1052631578947367 z"/>
                                <path fill="#9be9a8" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.1052631578947367 1.7,2.1052631578947367 z"/>
                            </g>
                            <g transform="translate(-8.5, 10.052631578947368)">
                                <path fill="#30a14e" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#30a14e" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.9473684210526314 0,1.9473684210526314 z"/>
                                <path fill="#30a14e" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.9473684210526314 1.7,2.9473684210526314 z"/>
                            </g>
                            <g transform="translate(-10.2, 12)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                        </g>
                        <g transform="translate(13.6, 8)">
                            <g transform="translate(0, 6)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-1.7, 6.2631578947368425)">
                                <path fill="#30a14e" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#30a14e" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.736842105263158 0,1.736842105263158 z"/>
                                <path fill="#30a14e" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.736842105263158 1.7,2.736842105263158 z"/>
                            </g>
                            <g transform="translate(-3.4, 7.473684210526315)">
                                <path fill="#40c463" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#40c463" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.526315789473684 0,1.526315789473684 z"/>
                                <path fill="#40c463" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.526315789473684 1.7,2.526315789473684 z"/>
                            </g>
                            <g transform="translate(-5.1, 8.368421052631579)">
                                <path fill="#40c463" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#40c463" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.6315789473684212 0,1.631578947368421 z"/>
                                <path fill="#40c463" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.631578947368421 1.7,2.6315789473684212 z"/>
                            </g>
                            <g transform="translate(-6.8, 9.578947368421053)">
                                <path fill="#40c463" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#40c463" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.4210526315789473 0,1.4210526315789473 z"/>
                                <path fill="#40c463" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.4210526315789473 1.7,2.4210526315789473 z"/>
                            </g>
                            <g transform="translate(-8.5, 11)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-10.2, 11.894736842105264)">
                                <path fill="#9be9a8" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#9be9a8" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.1052631578947367 0,1.1052631578947367 z"/>
                                <path fill="#9be9a8" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.1052631578947367 1.7,2.1052631578947367 z"/>
                            </g>
                        </g>
                        <g transform="translate(15.299999999999999, 9)">
                            <g transform="translate(0, 6)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-1.7, 6.368421052631579)">
                                <path fill="#40c463" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#40c463" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.6315789473684212 0,1.631578947368421 z"/>
                                <path fill="#40c463" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.631578947368421 1.7,2.6315789473684212 z"/>
                            </g>
                            <g transform="translate(-3.4, 7.578947368421053)">
                                <path fill="#40c463" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#40c463" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.4210526315789473 0,1.4210526315789473 z"/>
                                <path fill="#40c463" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.4210526315789473 1.7,2.4210526315789473 z"/>
                            </g>
                            <g transform="translate(-5.1, 7.947368421052632)">
                                <path fill="#216e39" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#216e39" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,3.052631578947368 0,2.052631578947368 z"/>
                                <path fill="#216e39" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,2.052631578947368 1.7,3.052631578947368 z"/>
                            </g>
                            <g transform="translate(-6.8, 9.157894736842106)">
                                <path fill="#30a14e" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#30a14e" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.8421052631578947 0,1.8421052631578947 z"/>
                                <path fill="#30a14e" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.8421052631578947 1.7,2.8421052631578947 z"/>
                            </g>
                            <g transform="translate(-8.5, 10.052631578947368)">
                                <path fill="#30a14e" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#30a14e" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.9473684210526314 0,1.9473684210526314 z"/>
                                <path fill="#30a14e" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.9473684210526314 1.7,2.9473684210526314 z"/>
                            </g>
                            <g transform="translate(-10.2, 11.578947368421053)">
                                <path fill="#40c463" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#40c463" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.4210526315789473 0,1.4210526315789473 z"/>
                                <path fill="#40c463" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.4210526315789473 1.7,2.4210526315789473 z"/>
                            </g>
                        </g>
                        <g transform="translate(17, 10)">
                            <g transform="translate(0, 5.894736842105263)">
                                <path fill="#9be9a8" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#9be9a8" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.1052631578947367 0,1.1052631578947367 z"/>
                                <path fill="#9be9a8" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.1052631578947367 1.7,2.1052631578947367 z"/>
                            </g>
                            <g transform="translate(-1.7, 6.473684210526315)">
                                <path fill="#40c463" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#40c463" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.526315789473684 0,1.526315789473684 z"/>
                                <path fill="#40c463" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.526315789473684 1.7,2.526315789473684 z"/>
                            </g>
                            <g transform="translate(-3.4, 7.894736842105263)">
                                <path fill="#9be9a8" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#9be9a8" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.1052631578947367 0,1.1052631578947367 z"/>
                                <path fill="#9be9a8" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.1052631578947367 1.7,2.1052631578947367 z"/>
                            </g>
                            <g transform="translate(-5.1, 8.473684210526315)">
                                <path fill="#40c463" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#40c463" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.526315789473684 0,1.526315789473684 z"/>
                                <path fill="#40c463" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.526315789473684 1.7,2.526315789473684 z"/>
                            </g>
                            <g transform="translate(-6.8, 9.789473684210527)">
                                <path fill="#9be9a8" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#9be9a8" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.2105263157894735 0,1.2105263157894737 z"/>
                                <path fill="#9be9a8" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.2105263157894737 1.7,2.2105263157894735 z"/>
                            </g>
                            <g transform="translate(-8.5, 10.263157894736842)">
                                <path fill="#30a14e" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#30a14e" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.736842105263158 0,1.736842105263158 z"/>
                                <path fill="#30a14e" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.736842105263158 1.7,2.736842105263158 z"/>
                            </g>
                            <g transform="translate(-10.2, 11.263157894736842)">
                                <path fill="#30a14e" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#30a14e" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.736842105263158 0,1.736842105263158 z"/>
                                <path fill="#30a14e" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.736842105263158 1.7,2.736842105263158 z"/>
                            </g>
                        </g>
                        <g transform="translate(18.7, 11)">
                            <g transform="translate(0, 6)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-1.7, 6.157894736842105)">
                                <path fill="#30a14e" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#30a14e" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.8421052631578947 0,1.8421052631578947 z"/>
                                <path fill="#30a14e" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.8421052631578947 1.7,2.8421052631578947 z"/>
                            </g>
                            <g transform="translate(-3.4, 6.631578947368421)">
                                <path fill="#216e39" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#216e39" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,3.3684210526315788 0,2.3684210526315788 z"/>
                                <path fill="#216e39" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,2.3684210526315788 1.7,3.3684210526315788 z"/>
                            </g>
                            <g transform="translate(-5.1, 8.68421052631579)">
                                <path fill="#9be9a8" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#9be9a8" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.3157894736842106 0,1.3157894736842106 z"/>
                                <path fill="#9be9a8" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.3157894736842106 1.7,2.3157894736842106 z"/>
                            </g>
                            <g transform="translate(-6.8, 9.894736842105264)">
                                <path fill="#9be9a8" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#9be9a8" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.1052631578947367 0,1.1052631578947367 z"/>
                                <path fill="#9be9a8" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.1052631578947367 1.7,2.1052631578947367 z"/>
                            </g>
                            <g transform="translate(-8.5, 11)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-10.2, 12)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                        </g>
                        <g transform="translate(20.4, 12)">
                            <g transform="translate(0, 6)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-1.7, 5.947368421052632)">
                                <path fill="#216e39" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#216e39" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,3.052631578947368 0,2.052631578947368 z"/>
                                <path fill="#216e39" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,2.052631578947368 1.7,3.052631578947368 z"/>
                            </g>
                            <g transform="translate(-3.4, 7.157894736842105)">
                                <path fill="#30a14e" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#30a14e" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.8421052631578947 0,1.8421052631578947 z"/>
                                <path fill="#30a14e" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.8421052631578947 1.7,2.8421052631578947 z"/>
                            </g>
                            <g transform="translate(-5.1, 7.947368421052632)">
                                <path fill="#216e39" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#216e39" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,3.052631578947368 0,2.052631578947368 z"/>
                                <path fill="#216e39" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,2.052631578947368 1.7,3.052631578947368 z"/>
                            </g>
                            <g transform="translate(-6.8, 9.157894736842106)">
                                <path fill="#30a14e" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#30a14e" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.8421052631578947 0,1.8421052631578947 z"/>
                                <path fill="#30a14e" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.8421052631578947 1.7,2.8421052631578947 z"/>
                            </g>
                            <g transform="translate(-8.5, 9.631578947368421)">
                                <path fill="#216e39" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#216e39" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,3.3684210526315788 0,2.3684210526315788 z"/>
                                <path fill="#216e39" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,2.3684210526315788 1.7,3.3684210526315788 z"/>
                            </g>
                            <g transform="translate(-10.2, 11.789473684210527)">
                                <path fill="#9be9a8" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#9be9a8" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.2105263157894735 0,1.2105263157894737 z"/>
                                <path fill="#9be9a8" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.2105263157894737 1.7,2.2105263157894735 z"/>
                            </g>
                        </g>
                        <g transform="translate(22.099999999999998, 13)">
                            <g transform="translate(0, 6)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-1.7, 7)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-3.4, 8)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-5.1, 9)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-6.8, 8.842105263157896)">
                                <path fill="#216e39" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#216e39" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,3.1578947368421053 0,2.1578947368421053 z"/>
                                <path fill="#216e39" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,2.1578947368421053 1.7,3.1578947368421053 z"/>
                            </g>
                            <g transform="translate(-8.5, 9.631578947368421)">
                                <path fill="#216e39" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#216e39" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,3.3684210526315788 0,2.3684210526315788 z"/>
                                <path fill="#216e39" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,2.3684210526315788 1.7,3.3684210526315788 z"/>
                            </g>
                            <g transform="translate(-10.2, 11.789473684210527)">
                                <path fill="#9be9a8" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#9be9a8" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.2105263157894735 0,1.2105263157894737 z"/>
                                <path fill="#9be9a8" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.2105263157894737 1.7,2.2105263157894735 z"/>
                            </g>
                        </g>
                        <g transform="translate(23.8, 14)">
                            <g transform="translate(0, 6)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-1.7, 5.842105263157896)">
                                <path fill="#216e39" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#216e39" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,3.1578947368421053 0,2.1578947368421053 z"/>
                                <path fill="#216e39" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,2.1578947368421053 1.7,3.1578947368421053 z"/>
                            </g>
                            <g transform="translate(-3.4, 8)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-5.1, 8.473684210526315)">
                                <path fill="#40c463" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#40c463" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.526315789473684 0,1.526315789473684 z"/>
                                <path fill="#40c463" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.526315789473684 1.7,2.526315789473684 z"/>
                            </g>
                            <g transform="translate(-6.8, 9.052631578947368)">
                                <path fill="#30a14e" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#30a14e" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.9473684210526314 0,1.9473684210526314 z"/>
                                <path fill="#30a14e" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.9473684210526314 1.7,2.9473684210526314 z"/>
                            </g>
                            <g transform="translate(-8.5, 10.578947368421053)">
                                <path fill="#40c463" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#40c463" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.4210526315789473 0,1.4210526315789473 z"/>
                                <path fill="#40c463" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.4210526315789473 1.7,2.4210526315789473 z"/>
                            </g>
                            <g transform="translate(-10.2, 12)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                        </g>
                        <g transform="translate(25.5, 15)">
                            <g transform="translate(0, 6)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-1.7, 6.052631578947368)">
                                <path fill="#30a14e" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#30a14e" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.9473684210526314 0,1.9473684210526314 z"/>
                                <path fill="#30a14e" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.9473684210526314 1.7,2.9473684210526314 z"/>
                            </g>
                            <g transform="translate(-3.4, 6.842105263157896)">
                                <path fill="#216e39" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#216e39" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,3.1578947368421053 0,2.1578947368421053 z"/>
                                <path fill="#216e39" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,2.1578947368421053 1.7,3.1578947368421053 z"/>
                            </g>
                            <g transform="translate(-5.1, 8.052631578947368)">
                                <path fill="#30a14e" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#30a14e" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.9473684210526314 0,1.9473684210526314 z"/>
                                <path fill="#30a14e" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.9473684210526314 1.7,2.9473684210526314 z"/>
                            </g>
                            <g transform="translate(-6.8, 9.68421052631579)">
                                <path fill="#9be9a8" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#9be9a8" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.3157894736842106 0,1.3157894736842106 z"/>
                                <path fill="#9be9a8" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.3157894736842106 1.7,2.3157894736842106 z"/>
                            </g>
                            <g transform="translate(-8.5, 10.578947368421053)">
                                <path fill="#40c463" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#40c463" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.4210526315789473 0,1.4210526315789473 z"/>
                                <path fill="#40c463" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.4210526315789473 1.7,2.4210526315789473 z"/>
                            </g>
                            <g transform="translate(-10.2, 11.68421052631579)">
                                <path fill="#9be9a8" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#9be9a8" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.3157894736842106 0,1.3157894736842106 z"/>
                                <path fill="#9be9a8" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.3157894736842106 1.7,2.3157894736842106 z"/>
                            </g>
                        </g>
                        <g transform="translate(27.2, 16)">
                            <g transform="translate(0, 5.578947368421053)">
                                <path fill="#9be9a8" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#9be9a8" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.4210526315789473 0,1.4210526315789473 z"/>
                                <path fill="#9be9a8" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.4210526315789473 1.7,2.4210526315789473 z"/>
                            </g>
                            <g transform="translate(-1.7, 6.473684210526315)">
                                <path fill="#40c463" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#40c463" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.526315789473684 0,1.526315789473684 z"/>
                                <path fill="#40c463" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.526315789473684 1.7,2.526315789473684 z"/>
                            </g>
                            <g transform="translate(-3.4, 6.7368421052631575)">
                                <path fill="#30a14e" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#30a14e" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,3.263157894736842 0,2.263157894736842 z"/>
                                <path fill="#30a14e" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,2.263157894736842 1.7,3.263157894736842 z"/>
                            </g>
                            <g transform="translate(-5.1, 8.263157894736842)">
                                <path fill="#40c463" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#40c463" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.736842105263158 0,1.736842105263158 z"/>
                                <path fill="#40c463" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.736842105263158 1.7,2.736842105263158 z"/>
                            </g>
                            <g transform="translate(-6.8, 9.473684210526315)">
                                <path fill="#40c463" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#40c463" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.526315789473684 0,1.526315789473684 z"/>
                                <path fill="#40c463" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.526315789473684 1.7,2.526315789473684 z"/>
                            </g>
                            <g transform="translate(-8.5, 10.263157894736842)">
                                <path fill="#40c463" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#40c463" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.736842105263158 0,1.736842105263158 z"/>
                                <path fill="#40c463" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.736842105263158 1.7,2.736842105263158 z"/>
                            </g>
                            <g transform="translate(-10.2, 12)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                        </g>
                        <g transform="translate(28.9, 17)">
                            <g transform="translate(0, 6)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-1.7, 6.052631578947368)">
                                <path fill="#30a14e" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#30a14e" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.9473684210526314 0,1.9473684210526314 z"/>
                                <path fill="#30a14e" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.9473684210526314 1.7,2.9473684210526314 z"/>
                            </g>
                            <g transform="translate(-3.4, 6.947368421052632)">
                                <path fill="#30a14e" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#30a14e" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,3.052631578947368 0,2.052631578947368 z"/>
                                <path fill="#30a14e" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,2.052631578947368 1.7,3.052631578947368 z"/>
                            </g>
                            <g transform="translate(-5.1, 7.947368421052632)">
                                <path fill="#30a14e" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#30a14e" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,3.052631578947368 0,2.052631578947368 z"/>
                                <path fill="#30a14e" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,2.052631578947368 1.7,3.052631578947368 z"/>
                            </g>
                            <g transform="translate(-6.8, 9.052631578947368)">
                                <path fill="#30a14e" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#30a14e" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.9473684210526314 0,1.9473684210526314 z"/>
                                <path fill="#30a14e" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.9473684210526314 1.7,2.9473684210526314 z"/>
                            </g>
                            <g transform="translate(-8.5, 9.210526315789473)">
                                <path fill="#216e39" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#216e39" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,3.789473684210526 0,2.789473684210526 z"/>
                                <path fill="#216e39" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,2.789473684210526 1.7,3.789473684210526 z"/>
                            </g>
                            <g transform="translate(-10.2, 12)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                        </g>
                        <g transform="translate(30.599999999999998, 18)">
                            <g transform="translate(0, 5.684210526315789)">
                                <path fill="#9be9a8" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#9be9a8" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.3157894736842106 0,1.3157894736842106 z"/>
                                <path fill="#9be9a8" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.3157894736842106 1.7,2.3157894736842106 z"/>
                            </g>
                            <g transform="translate(-1.7, 7)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-3.4, 6.947368421052632)">
                                <path fill="#30a14e" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#30a14e" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,3.052631578947368 0,2.052631578947368 z"/>
                                <path fill="#30a14e" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,2.052631578947368 1.7,3.052631578947368 z"/>
                            </g>
                            <g transform="translate(-5.1, 8.578947368421053)">
                                <path fill="#9be9a8" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#9be9a8" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.4210526315789473 0,1.4210526315789473 z"/>
                                <path fill="#9be9a8" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.4210526315789473 1.7,2.4210526315789473 z"/>
                            </g>
                            <g transform="translate(-6.8, 8.947368421052632)">
                                <path fill="#30a14e" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#30a14e" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,3.052631578947368 0,2.052631578947368 z"/>
                                <path fill="#30a14e" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,2.052631578947368 1.7,3.052631578947368 z"/>
                            </g>
                            <g transform="translate(-8.5, 10.68421052631579)">
                                <path fill="#9be9a8" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#9be9a8" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.3157894736842106 0,1.3157894736842106 z"/>
                                <path fill="#9be9a8" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.3157894736842106 1.7,2.3157894736842106 z"/>
                            </g>
                            <g transform="translate(-10.2, 10.526315789473685)">
                                <path fill="#216e39" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#216e39" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,3.473684210526316 0,2.473684210526316 z"/>
                                <path fill="#216e39" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,2.473684210526316 1.7,3.473684210526316 z"/>
                            </g>
                        </g>
                        <g transform="translate(32.3, 19)">
                            <g transform="translate(0, 5.052631578947368)">
                                <path fill="#30a14e" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#30a14e" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.9473684210526314 0,1.9473684210526314 z"/>
                                <path fill="#30a14e" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.9473684210526314 1.7,2.9473684210526314 z"/>
                            </g>
                            <g transform="translate(-1.7, 6.2631578947368425)">
                                <path fill="#40c463" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#40c463" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.736842105263158 0,1.736842105263158 z"/>
                                <path fill="#40c463" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.736842105263158 1.7,2.736842105263158 z"/>
                            </g>
                            <g transform="translate(-3.4, 6.947368421052632)">
                                <path fill="#30a14e" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#30a14e" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,3.052631578947368 0,2.052631578947368 z"/>
                                <path fill="#30a14e" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,2.052631578947368 1.7,3.052631578947368 z"/>
                            </g>
                            <g transform="translate(-5.1, 8.052631578947368)">
                                <path fill="#30a14e" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#30a14e" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.9473684210526314 0,1.9473684210526314 z"/>
                                <path fill="#30a14e" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.9473684210526314 1.7,2.9473684210526314 z"/>
                            </g>
                            <g transform="translate(-6.8, 9.894736842105264)">
                                <path fill="#9be9a8" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#9be9a8" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.1052631578947367 0,1.1052631578947367 z"/>
                                <path fill="#9be9a8" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.1052631578947367 1.7,2.1052631578947367 z"/>
                            </g>
                            <g transform="translate(-8.5, 10.894736842105264)">
                                <path fill="#9be9a8" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#9be9a8" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.1052631578947367 0,1.1052631578947367 z"/>
                                <path fill="#9be9a8" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.1052631578947367 1.7,2.1052631578947367 z"/>
                            </g>
                            <g transform="translate(-10.2, 12)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                        </g>
                        <g transform="translate(34, 20)">
                            <g transform="translate(0, 5.894736842105263)">
                                <path fill="#9be9a8" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#9be9a8" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.1052631578947367 0,1.1052631578947367 z"/>
                                <path fill="#9be9a8" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.1052631578947367 1.7,2.1052631578947367 z"/>
                            </g>
                            <g transform="translate(-1.7, 5.526315789473684)">
                                <path fill="#216e39" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#216e39" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,3.473684210526316 0,2.473684210526316 z"/>
                                <path fill="#216e39" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,2.473684210526316 1.7,3.473684210526316 z"/>
                            </g>
                            <g transform="translate(-3.4, 6.7368421052631575)">
                                <path fill="#30a14e" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#30a14e" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,3.263157894736842 0,2.263157894736842 z"/>
                                <path fill="#30a14e" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,2.263157894736842 1.7,3.263157894736842 z"/>
                            </g>
                            <g transform="translate(-5.1, 7.7368421052631575)">
                                <path fill="#30a14e" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#30a14e" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,3.263157894736842 0,2.263157894736842 z"/>
                                <path fill="#30a14e" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,2.263157894736842 1.7,3.263157894736842 z"/>
                            </g>
                            <g transform="translate(-6.8, 9.68421052631579)">
                                <path fill="#9be9a8" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#9be9a8" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.3157894736842106 0,1.3157894736842106 z"/>
                                <path fill="#9be9a8" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.3157894736842106 1.7,2.3157894736842106 z"/>
                            </g>
                            <g transform="translate(-8.5, 10.578947368421053)">
                                <path fill="#9be9a8" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#9be9a8" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.4210526315789473 0,1.4210526315789473 z"/>
                                <path fill="#9be9a8" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.4210526315789473 1.7,2.4210526315789473 z"/>
                            </g>
                            <g transform="translate(-10.2, 11.894736842105264)">
                                <path fill="#9be9a8" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#9be9a8" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.1052631578947367 0,1.1052631578947367 z"/>
                                <path fill="#9be9a8" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.1052631578947367 1.7,2.1052631578947367 z"/>
                            </g>
                        </g>
                        <g transform="translate(35.699999999999996, 21)">
                            <g transform="translate(0, 6)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-1.7, 6.052631578947368)">
                                <path fill="#30a14e" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#30a14e" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.9473684210526314 0,1.9473684210526314 z"/>
                                <path fill="#30a14e" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.9473684210526314 1.7,2.9473684210526314 z"/>
                            </g>
                            <g transform="translate(-3.4, 6.947368421052632)">
                                <path fill="#30a14e" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#30a14e" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,3.052631578947368 0,2.052631578947368 z"/>
                                <path fill="#30a14e" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,2.052631578947368 1.7,3.052631578947368 z"/>
                            </g>
                            <g transform="translate(-5.1, 9)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-6.8, 9.578947368421053)">
                                <path fill="#9be9a8" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#9be9a8" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.4210526315789473 0,1.4210526315789473 z"/>
                                <path fill="#9be9a8" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.4210526315789473 1.7,2.4210526315789473 z"/>
                            </g>
                            <g transform="translate(-8.5, 10.578947368421053)">
                                <path fill="#9be9a8" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#9be9a8" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.4210526315789473 0,1.4210526315789473 z"/>
                                <path fill="#9be9a8" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.4210526315789473 1.7,2.4210526315789473 z"/>
                            </g>
                            <g transform="translate(-10.2, 11.894736842105264)">
                                <path fill="#9be9a8" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#9be9a8" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.1052631578947367 0,1.1052631578947367 z"/>
                                <path fill="#9be9a8" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.1052631578947367 1.7,2.1052631578947367 z"/>
                            </g>
                        </g>
                        <g transform="translate(37.4, 22)">
                            <g transform="translate(0, 5.684210526315789)">
                                <path fill="#9be9a8" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#9be9a8" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.3157894736842106 0,1.3157894736842106 z"/>
                                <path fill="#9be9a8" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.3157894736842106 1.7,2.3157894736842106 z"/>
                            </g>
                            <g transform="translate(-1.7, 6.684210526315789)">
                                <path fill="#9be9a8" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#9be9a8" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.3157894736842106 0,1.3157894736842106 z"/>
                                <path fill="#9be9a8" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.3157894736842106 1.7,2.3157894736842106 z"/>
                            </g>
                            <g transform="translate(-3.4, 7.7894736842105265)">
                                <path fill="#9be9a8" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#9be9a8" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.2105263157894735 0,1.2105263157894737 z"/>
                                <path fill="#9be9a8" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.2105263157894737 1.7,2.2105263157894735 z"/>
                            </g>
                            <g transform="translate(-5.1, 8.578947368421053)">
                                <path fill="#9be9a8" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#9be9a8" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.4210526315789473 0,1.4210526315789473 z"/>
                                <path fill="#9be9a8" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.4210526315789473 1.7,2.4210526315789473 z"/>
                            </g>
                            <g transform="translate(-6.8, 9.368421052631579)">
                                <path fill="#40c463" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#40c463" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.6315789473684212 0,1.631578947368421 z"/>
                                <path fill="#40c463" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.631578947368421 1.7,2.6315789473684212 z"/>
                            </g>
                            <g transform="translate(-8.5, 11)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-10.2, 12)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                        </g>
                        <g transform="translate(39.1, 23)">
                            <g transform="translate(0, 6)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-1.7, 5.7368421052631575)">
                                <path fill="#30a14e" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#30a14e" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,3.263157894736842 0,2.263157894736842 z"/>
                                <path fill="#30a14e" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,2.263157894736842 1.7,3.263157894736842 z"/>
                            </g>
                            <g transform="translate(-3.4, 7.684210526315789)">
                                <path fill="#9be9a8" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#9be9a8" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.3157894736842106 0,1.3157894736842106 z"/>
                                <path fill="#9be9a8" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.3157894736842106 1.7,2.3157894736842106 z"/>
                            </g>
                            <g transform="translate(-5.1, 8.157894736842106)">
                                <path fill="#40c463" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#40c463" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.8421052631578947 0,1.8421052631578947 z"/>
                                <path fill="#40c463" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.8421052631578947 1.7,2.8421052631578947 z"/>
                            </g>
                            <g transform="translate(-6.8, 8.947368421052632)">
                                <path fill="#30a14e" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#30a14e" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,3.052631578947368 0,2.052631578947368 z"/>
                                <path fill="#30a14e" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,2.052631578947368 1.7,3.052631578947368 z"/>
                            </g>
                            <g transform="translate(-8.5, 9.210526315789473)">
                                <path fill="#216e39" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#216e39" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,3.789473684210526 0,2.789473684210526 z"/>
                                <path fill="#216e39" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,2.789473684210526 1.7,3.789473684210526 z"/>
                            </g>
                            <g transform="translate(-10.2, 12)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                        </g>
                        <g transform="translate(40.8, 24)">
                            <g transform="translate(0, 6)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-1.7, 6.052631578947368)">
                                <path fill="#30a14e" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#30a14e" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.9473684210526314 0,1.9473684210526314 z"/>
                                <path fill="#30a14e" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.9473684210526314 1.7,2.9473684210526314 z"/>
                            </g>
                            <g transform="translate(-3.4, 7.2631578947368425)">
                                <path fill="#40c463" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#40c463" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.736842105263158 0,1.736842105263158 z"/>
                                <path fill="#40c463" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.736842105263158 1.7,2.736842105263158 z"/>
                            </g>
                            <g transform="translate(-5.1, 7.842105263157896)">
                                <path fill="#30a14e" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#30a14e" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,3.1578947368421053 0,2.1578947368421053 z"/>
                                <path fill="#30a14e" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,2.1578947368421053 1.7,3.1578947368421053 z"/>
                            </g>
                            <g transform="translate(-6.8, 8.210526315789473)">
                                <path fill="#216e39" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#216e39" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,3.789473684210526 0,2.789473684210526 z"/>
                                <path fill="#216e39" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,2.789473684210526 1.7,3.789473684210526 z"/>
                            </g>
                            <g transform="translate(-8.5, 10.157894736842106)">
                                <path fill="#40c463" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#40c463" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.8421052631578947 0,1.8421052631578947 z"/>
                                <path fill="#40c463" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.8421052631578947 1.7,2.8421052631578947 z"/>
                            </g>
                            <g transform="translate(-10.2, 11.894736842105264)">
                                <path fill="#9be9a8" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#9be9a8" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.1052631578947367 0,1.1052631578947367 z"/>
                                <path fill="#9be9a8" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.1052631578947367 1.7,2.1052631578947367 z"/>
                            </g>
                        </g>
                        <g transform="translate(42.5, 25)">
                            <g transform="translate(0, 6)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-1.7, 6.578947368421053)">
                                <path fill="#9be9a8" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#9be9a8" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.4210526315789473 0,1.4210526315789473 z"/>
                                <path fill="#9be9a8" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.4210526315789473 1.7,2.4210526315789473 z"/>
                            </g>
                            <g transform="translate(-3.4, 6.842105263157896)">
                                <path fill="#30a14e" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#30a14e" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,3.1578947368421053 0,2.1578947368421053 z"/>
                                <path fill="#30a14e" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,2.1578947368421053 1.7,3.1578947368421053 z"/>
                            </g>
                            <g transform="translate(-5.1, 7.842105263157896)">
                                <path fill="#30a14e" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#30a14e" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,3.1578947368421053 0,2.1578947368421053 z"/>
                                <path fill="#30a14e" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,2.1578947368421053 1.7,3.1578947368421053 z"/>
                            </g>
                            <g transform="translate(-6.8, 9.68421052631579)">
                                <path fill="#9be9a8" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#9be9a8" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.3157894736842106 0,1.3157894736842106 z"/>
                                <path fill="#9be9a8" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.3157894736842106 1.7,2.3157894736842106 z"/>
                            </g>
                            <g transform="translate(-8.5, 9.421052631578949)">
                                <path fill="#216e39" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#216e39" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,3.5789473684210527 0,2.5789473684210527 z"/>
                                <path fill="#216e39" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,2.5789473684210527 1.7,3.5789473684210527 z"/>
                            </g>
                            <g transform="translate(-10.2, 12)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                        </g>
                        <g transform="translate(44.199999999999996, 26)">
                            <g transform="translate(0, 5.578947368421053)">
                                <path fill="#9be9a8" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#9be9a8" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.4210526315789473 0,1.4210526315789473 z"/>
                                <path fill="#9be9a8" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.4210526315789473 1.7,2.4210526315789473 z"/>
                            </g>
                            <g transform="translate(-1.7, 5.947368421052632)">
                                <path fill="#30a14e" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#30a14e" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,3.052631578947368 0,2.052631578947368 z"/>
                                <path fill="#30a14e" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,2.052631578947368 1.7,3.052631578947368 z"/>
                            </g>
                            <g transform="translate(-3.4, 7.2631578947368425)">
                                <path fill="#40c463" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#40c463" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.736842105263158 0,1.736842105263158 z"/>
                                <path fill="#40c463" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.736842105263158 1.7,2.736842105263158 z"/>
                            </g>
                            <g transform="translate(-5.1, 8.368421052631579)">
                                <path fill="#40c463" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#40c463" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.6315789473684212 0,1.631578947368421 z"/>
                                <path fill="#40c463" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.631578947368421 1.7,2.6315789473684212 z"/>
                            </g>
                            <g transform="translate(-6.8, 9.263157894736842)">
                                <path fill="#40c463" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#40c463" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.736842105263158 0,1.736842105263158 z"/>
                                <path fill="#40c463" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.736842105263158 1.7,2.736842105263158 z"/>
                            </g>
                            <g transform="translate(-8.5, 11)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-10.2, 12)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                        </g>
                        <g transform="translate(45.9, 27)">
                            <g transform="translate(0, 5.894736842105263)">
                                <path fill="#9be9a8" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#9be9a8" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.1052631578947367 0,1.1052631578947367 z"/>
                                <path fill="#9be9a8" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.1052631578947367 1.7,2.1052631578947367 z"/>
                            </g>
                            <g transform="translate(-1.7, 6.684210526315789)">
                                <path fill="#9be9a8" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#9be9a8" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.3157894736842106 0,1.3157894736842106 z"/>
                                <path fill="#9be9a8" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.3157894736842106 1.7,2.3157894736842106 z"/>
                            </g>
                            <g transform="translate(-3.4, 7.684210526315789)">
                                <path fill="#9be9a8" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#9be9a8" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.3157894736842106 0,1.3157894736842106 z"/>
                                <path fill="#9be9a8" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.3157894736842106 1.7,2.3157894736842106 z"/>
                            </g>
                            <g transform="translate(-5.1, 8.052631578947368)">
                                <path fill="#30a14e" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#30a14e" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.9473684210526314 0,1.9473684210526314 z"/>
                                <path fill="#30a14e" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.9473684210526314 1.7,2.9473684210526314 z"/>
                            </g>
                            <g transform="translate(-6.8, 9.68421052631579)">
                                <path fill="#9be9a8" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#9be9a8" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.3157894736842106 0,1.3157894736842106 z"/>
                                <path fill="#9be9a8" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.3157894736842106 1.7,2.3157894736842106 z"/>
                            </g>
                            <g transform="translate(-8.5, 10.68421052631579)">
                                <path fill="#9be9a8" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#9be9a8" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.3157894736842106 0,1.3157894736842106 z"/>
                                <path fill="#9be9a8" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.3157894736842106 1.7,2.3157894736842106 z"/>
                            </g>
                            <g transform="translate(-10.2, 12)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                        </g>
                        <g transform="translate(47.6, 28)">
                            <g transform="translate(0, 6)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-1.7, 5.7368421052631575)">
                                <path fill="#216e39" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#216e39" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,3.263157894736842 0,2.263157894736842 z"/>
                                <path fill="#216e39" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,2.263157894736842 1.7,3.263157894736842 z"/>
                            </g>
                            <g transform="translate(-3.4, 7.7894736842105265)">
                                <path fill="#9be9a8" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#9be9a8" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.2105263157894735 0,1.2105263157894737 z"/>
                                <path fill="#9be9a8" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.2105263157894737 1.7,2.2105263157894735 z"/>
                            </g>
                            <g transform="translate(-5.1, 8.052631578947368)">
                                <path fill="#30a14e" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#30a14e" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.9473684210526314 0,1.9473684210526314 z"/>
                                <path fill="#30a14e" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.9473684210526314 1.7,2.9473684210526314 z"/>
                            </g>
                            <g transform="translate(-6.8, 9.789473684210527)">
                                <path fill="#9be9a8" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#9be9a8" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.2105263157894735 0,1.2105263157894737 z"/>
                                <path fill="#9be9a8" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.2105263157894737 1.7,2.2105263157894735 z"/>
                            </g>
                            <g transform="translate(-8.5, 10.368421052631579)">
                                <path fill="#40c463" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#40c463" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.6315789473684212 0,1.631578947368421 z"/>
                                <path fill="#40c463" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.631578947368421 1.7,2.6315789473684212 z"/>
                            </g>
                            <g transform="translate(-10.2, 11.894736842105264)">
                                <path fill="#9be9a8" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#9be9a8" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.1052631578947367 0,1.1052631578947367 z"/>
                                <path fill="#9be9a8" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.1052631578947367 1.7,2.1052631578947367 z"/>
                            </g>
                        </g>
                        <g transform="translate(49.3, 29)">
                            <g transform="translate(0, 6)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-1.7, 6.7894736842105265)">
                                <path fill="#9be9a8" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#9be9a8" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.2105263157894735 0,1.2105263157894737 z"/>
                                <path fill="#9be9a8" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.2105263157894737 1.7,2.2105263157894735 z"/>
                            </g>
                            <g transform="translate(-3.4, 7.7894736842105265)">
                                <path fill="#9be9a8" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#9be9a8" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.2105263157894735 0,1.2105263157894737 z"/>
                                <path fill="#9be9a8" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.2105263157894737 1.7,2.2105263157894735 z"/>
                            </g>
                            <g transform="translate(-5.1, 8.052631578947368)">
                                <path fill="#30a14e" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#30a14e" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.9473684210526314 0,1.9473684210526314 z"/>
                                <path fill="#30a14e" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.9473684210526314 1.7,2.9473684210526314 z"/>
                            </g>
                            <g transform="translate(-6.8, 9.157894736842106)">
                                <path fill="#30a14e" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#30a14e" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.8421052631578947 0,1.8421052631578947 z"/>
                                <path fill="#30a14e" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.8421052631578947 1.7,2.8421052631578947 z"/>
                            </g>
                            <g transform="translate(-8.5, 10.789473684210527)">
                                <path fill="#9be9a8" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#9be9a8" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.2105263157894735 0,1.2105263157894737 z"/>
                                <path fill="#9be9a8" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.2105263157894737 1.7,2.2105263157894735 z"/>
                            </g>
                            <g transform="translate(-10.2, 12)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                        </g>
                        <g transform="translate(51, 30)">
                            <g transform="translate(0, 5.894736842105263)">
                                <path fill="#9be9a8" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#9be9a8" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.1052631578947367 0,1.1052631578947367 z"/>
                                <path fill="#9be9a8" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.1052631578947367 1.7,2.1052631578947367 z"/>
                            </g>
                            <g transform="translate(-1.7, 6.052631578947368)">
                                <path fill="#30a14e" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#30a14e" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.9473684210526314 0,1.9473684210526314 z"/>
                                <path fill="#30a14e" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.9473684210526314 1.7,2.9473684210526314 z"/>
                            </g>
                            <g transform="translate(-3.4, 6.842105263157896)">
                                <path fill="#216e39" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#216e39" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,3.1578947368421053 0,2.1578947368421053 z"/>
                                <path fill="#216e39" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,2.1578947368421053 1.7,3.1578947368421053 z"/>
                            </g>
                            <g transform="translate(-5.1, 7.526315789473684)">
                                <path fill="#216e39" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#216e39" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,3.473684210526316 0,2.473684210526316 z"/>
                                <path fill="#216e39" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,2.473684210526316 1.7,3.473684210526316 z"/>
                            </g>
                            <g transform="translate(-6.8, 8.736842105263158)">
                                <path fill="#216e39" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#216e39" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,3.263157894736842 0,2.263157894736842 z"/>
                                <path fill="#216e39" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,2.263157894736842 1.7,3.263157894736842 z"/>
                            </g>
                            <g transform="translate(-8.5, 11)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-10.2, 12)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                        </g>
                        <g transform="translate(52.699999999999996, 31)">
                            <g transform="translate(0, 6)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-1.7, 7)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-3.4, 7.052631578947368)">
                                <path fill="#30a14e" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#30a14e" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.9473684210526314 0,1.9473684210526314 z"/>
                                <path fill="#30a14e" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.9473684210526314 1.7,2.9473684210526314 z"/>
                            </g>
                            <g transform="translate(-5.1, 8.368421052631579)">
                                <path fill="#40c463" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#40c463" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.6315789473684212 0,1.631578947368421 z"/>
                                <path fill="#40c463" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.631578947368421 1.7,2.6315789473684212 z"/>
                            </g>
                            <g transform="translate(-6.8, 8.736842105263158)">
                                <path fill="#216e39" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#216e39" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,3.263157894736842 0,2.263157894736842 z"/>
                                <path fill="#216e39" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,2.263157894736842 1.7,3.263157894736842 z"/>
                            </g>
                            <g transform="translate(-8.5, 10.157894736842106)">
                                <path fill="#30a14e" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#30a14e" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.8421052631578947 0,1.8421052631578947 z"/>
                                <path fill="#30a14e" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.8421052631578947 1.7,2.8421052631578947 z"/>
                            </g>
                            <g transform="translate(-10.2, 11.68421052631579)">
                                <path fill="#9be9a8" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#9be9a8" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.3157894736842106 0,1.3157894736842106 z"/>
                                <path fill="#9be9a8" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.3157894736842106 1.7,2.3157894736842106 z"/>
                            </g>
                        </g>
                        <g transform="translate(54.4, 32)">
                            <g transform="translate(0, 6)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-1.7, 6.578947368421053)">
                                <path fill="#9be9a8" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#9be9a8" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.4210526315789473 0,1.4210526315789473 z"/>
                                <path fill="#9be9a8" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.4210526315789473 1.7,2.4210526315789473 z"/>
                            </g>
                            <g transform="translate(-3.4, 7.473684210526315)">
                                <path fill="#40c463" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#40c463" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.526315789473684 0,1.526315789473684 z"/>
                                <path fill="#40c463" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.526315789473684 1.7,2.526315789473684 z"/>
                            </g>
                            <g transform="translate(-5.1, 8.68421052631579)">
                                <path fill="#9be9a8" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#9be9a8" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.3157894736842106 0,1.3157894736842106 z"/>
                                <path fill="#9be9a8" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.3157894736842106 1.7,2.3157894736842106 z"/>
                            </g>
                            <g transform="translate(-6.8, 8.842105263157896)">
                                <path fill="#30a14e" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#30a14e" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,3.1578947368421053 0,2.1578947368421053 z"/>
                                <path fill="#30a14e" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,2.1578947368421053 1.7,3.1578947368421053 z"/>
                            </g>
                            <g transform="translate(-8.5, 10.789473684210527)">
                                <path fill="#9be9a8" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#9be9a8" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.2105263157894735 0,1.2105263157894737 z"/>
                                <path fill="#9be9a8" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.2105263157894737 1.7,2.2105263157894735 z"/>
                            </g>
                            <g transform="translate(-10.2, 12)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                        </g>
                        <g transform="translate(56.1, 33)">
                            <g transform="translate(0, 6)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-1.7, 6.368421052631579)">
                                <path fill="#40c463" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#40c463" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.6315789473684212 0,1.631578947368421 z"/>
                                <path fill="#40c463" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.631578947368421 1.7,2.6315789473684212 z"/>
                            </g>
                            <g transform="translate(-3.4, 6.842105263157896)">
                                <path fill="#30a14e" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#30a14e" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,3.1578947368421053 0,2.1578947368421053 z"/>
                                <path fill="#30a14e" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,2.1578947368421053 1.7,3.1578947368421053 z"/>
                            </g>
                            <g transform="translate(-5.1, 8.578947368421053)">
                                <path fill="#9be9a8" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#9be9a8" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.4210526315789473 0,1.4210526315789473 z"/>
                                <path fill="#9be9a8" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.4210526315789473 1.7,2.4210526315789473 z"/>
                            </g>
                            <g transform="translate(-6.8, 9.473684210526315)">
                                <path fill="#40c463" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#40c463" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.526315789473684 0,1.526315789473684 z"/>
                                <path fill="#40c463" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.526315789473684 1.7,2.526315789473684 z"/>
                            </g>
                            <g transform="translate(-8.5, 10.473684210526315)">
                                <path fill="#40c463" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#40c463" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.526315789473684 0,1.526315789473684 z"/>
                                <path fill="#40c463" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.526315789473684 1.7,2.526315789473684 z"/>
                            </g>
                            <g transform="translate(-10.2, 11.68421052631579)">
                                <path fill="#9be9a8" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#9be9a8" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.3157894736842106 0,1.3157894736842106 z"/>
                                <path fill="#9be9a8" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.3157894736842106 1.7,2.3157894736842106 z"/>
                            </g>
                        </g>
                        <g transform="translate(57.8, 34)">
                            <g transform="translate(0, 5.684210526315789)">
                                <path fill="#9be9a8" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#9be9a8" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.3157894736842106 0,1.3157894736842106 z"/>
                                <path fill="#9be9a8" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.3157894736842106 1.7,2.3157894736842106 z"/>
                            </g>
                            <g transform="translate(-1.7, 5.105263157894737)">
                                <path fill="#216e39" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#216e39" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,3.894736842105263 0,2.894736842105263 z"/>
                                <path fill="#216e39" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,2.894736842105263 1.7,3.894736842105263 z"/>
                            </g>
                            <g transform="translate(-3.4, 7.157894736842105)">
                                <path fill="#40c463" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#40c463" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.8421052631578947 0,1.8421052631578947 z"/>
                                <path fill="#40c463" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.8421052631578947 1.7,2.8421052631578947 z"/>
                            </g>
                            <g transform="translate(-5.1, 9)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-6.8, 10)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-8.5, 11)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-10.2, 12)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                        </g>
                        <g transform="translate(59.5, 35)">
                            <g transform="translate(0, 6)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-1.7, 7)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-3.4, 7.684210526315789)">
                                <path fill="#9be9a8" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#9be9a8" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.3157894736842106 0,1.3157894736842106 z"/>
                                <path fill="#9be9a8" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.3157894736842106 1.7,2.3157894736842106 z"/>
                            </g>
                            <g transform="translate(-5.1, 7.526315789473684)">
                                <path fill="#216e39" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#216e39" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,3.473684210526316 0,2.473684210526316 z"/>
                                <path fill="#216e39" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,2.473684210526316 1.7,3.473684210526316 z"/>
                            </g>
                            <g transform="translate(-6.8, 9.368421052631579)">
                                <path fill="#40c463" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#40c463" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.6315789473684212 0,1.631578947368421 z"/>
                                <path fill="#40c463" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.631578947368421 1.7,2.6315789473684212 z"/>
                            </g>
                            <g transform="translate(-8.5, 10.263157894736842)">
                                <path fill="#40c463" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#40c463" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.736842105263158 0,1.736842105263158 z"/>
                                <path fill="#40c463" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.736842105263158 1.7,2.736842105263158 z"/>
                            </g>
                            <g transform="translate(-10.2, 11.578947368421053)">
                                <path fill="#9be9a8" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#9be9a8" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.4210526315789473 0,1.4210526315789473 z"/>
                                <path fill="#9be9a8" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.4210526315789473 1.7,2.4210526315789473 z"/>
                            </g>
                        </g>
                        <g transform="translate(61.199999999999996, 36)">
                            <g transform="translate(0, 6)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-1.7, 6.473684210526315)">
                                <path fill="#9be9a8" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#9be9a8" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.526315789473684 0,1.526315789473684 z"/>
                                <path fill="#9be9a8" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.526315789473684 1.7,2.526315789473684 z"/>
                            </g>
                            <g transform="translate(-3.4, 6)">
                                <path fill="#216e39" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#216e39" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,4 0,3 z"/>
                                <path fill="#216e39" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,3 1.7,4 z"/>
                            </g>
                            <g transform="translate(-5.1, 7.947368421052632)">
                                <path fill="#40c463" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#40c463" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,3.052631578947368 0,2.052631578947368 z"/>
                                <path fill="#40c463" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,2.052631578947368 1.7,3.052631578947368 z"/>
                            </g>
                            <g transform="translate(-6.8, 9.157894736842106)">
                                <path fill="#40c463" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#40c463" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.8421052631578947 0,1.8421052631578947 z"/>
                                <path fill="#40c463" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.8421052631578947 1.7,2.8421052631578947 z"/>
                            </g>
                            <g transform="translate(-8.5, 10.368421052631579)">
                                <path fill="#40c463" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#40c463" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.6315789473684212 0,1.631578947368421 z"/>
                                <path fill="#40c463" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.631578947368421 1.7,2.6315789473684212 z"/>
                            </g>
                            <g transform="translate(-10.2, 11.894736842105264)">
                                <path fill="#9be9a8" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#9be9a8" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.1052631578947367 0,1.1052631578947367 z"/>
                                <path fill="#9be9a8" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.1052631578947367 1.7,2.1052631578947367 z"/>
                            </g>
                        </g>
                        <g transform="translate(62.9, 37)">
                            <g transform="translate(0, 5.7894736842105265)">
                                <path fill="#9be9a8" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#9be9a8" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.2105263157894735 0,1.2105263157894737 z"/>
                                <path fill="#9be9a8" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.2105263157894737 1.7,2.2105263157894735 z"/>
                            </g>
                            <g transform="translate(-1.7, 6.157894736842105)">
                                <path fill="#40c463" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#40c463" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.8421052631578947 0,1.8421052631578947 z"/>
                                <path fill="#40c463" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.8421052631578947 1.7,2.8421052631578947 z"/>
                            </g>
                            <g transform="translate(-3.4, 7.2631578947368425)">
                                <path fill="#40c463" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#40c463" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.736842105263158 0,1.736842105263158 z"/>
                                <path fill="#40c463" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.736842105263158 1.7,2.736842105263158 z"/>
                            </g>
                            <g transform="translate(-5.1, 8.368421052631579)">
                                <path fill="#40c463" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#40c463" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.6315789473684212 0,1.631578947368421 z"/>
                                <path fill="#40c463" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.631578947368421 1.7,2.6315789473684212 z"/>
                            </g>
                            <g transform="translate(-6.8, 8.526315789473685)">
                                <path fill="#30a14e" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#30a14e" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,3.473684210526316 0,2.473684210526316 z"/>
                                <path fill="#30a14e" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,2.473684210526316 1.7,3.473684210526316 z"/>
                            </g>
                            <g transform="translate(-8.5, 9.31578947368421)">
                                <path fill="#216e39" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#216e39" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,3.6842105263157894 0,2.6842105263157894 z"/>
                                <path fill="#216e39" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,2.6842105263157894 1.7,3.6842105263157894 z"/>
                            </g>
                            <g transform="translate(-10.2, 11.68421052631579)">
                                <path fill="#9be9a8" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#9be9a8" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.3157894736842106 0,1.3157894736842106 z"/>
                                <path fill="#9be9a8" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.3157894736842106 1.7,2.3157894736842106 z"/>
                            </g>
                        </g>
                        <g transform="translate(64.6, 38)">
                            <g transform="translate(0, 5.368421052631579)">
                                <path fill="#40c463" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#40c463" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.6315789473684212 0,1.631578947368421 z"/>
                                <path fill="#40c463" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.631578947368421 1.7,2.6315789473684212 z"/>
                            </g>
                            <g transform="translate(-1.7, 6.7894736842105265)">
                                <path fill="#9be9a8" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#9be9a8" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.2105263157894735 0,1.2105263157894737 z"/>
                                <path fill="#9be9a8" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.2105263157894737 1.7,2.2105263157894735 z"/>
                            </g>
                            <g transform="translate(-3.4, 7.157894736842105)">
                                <path fill="#40c463" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#40c463" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.8421052631578947 0,1.8421052631578947 z"/>
                                <path fill="#40c463" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.8421052631578947 1.7,2.8421052631578947 z"/>
                            </g>
                            <g transform="translate(-5.1, 6.894736842105264)">
                                <path fill="#216e39" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#216e39" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,4.105263157894736 0,3.1052631578947367 z"/>
                                <path fill="#216e39" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,3.1052631578947367 1.7,4.105263157894736 z"/>
                            </g>
                            <g transform="translate(-6.8, 9.789473684210527)">
                                <path fill="#9be9a8" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#9be9a8" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.2105263157894735 0,1.2105263157894737 z"/>
                                <path fill="#9be9a8" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.2105263157894737 1.7,2.2105263157894735 z"/>
                            </g>
                            <g transform="translate(-8.5, 10.157894736842106)">
                                <path fill="#40c463" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#40c463" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.8421052631578947 0,1.8421052631578947 z"/>
                                <path fill="#40c463" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.8421052631578947 1.7,2.8421052631578947 z"/>
                            </g>
                            <g transform="translate(-10.2, 11.894736842105264)">
                                <path fill="#9be9a8" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#9be9a8" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.1052631578947367 0,1.1052631578947367 z"/>
                                <path fill="#9be9a8" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.1052631578947367 1.7,2.1052631578947367 z"/>
                            </g>
                        </g>
                        <g transform="translate(66.3, 39)">
                            <g transform="translate(0, 5.894736842105263)">
                                <path fill="#9be9a8" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#9be9a8" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.1052631578947367 0,1.1052631578947367 z"/>
                                <path fill="#9be9a8" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.1052631578947367 1.7,2.1052631578947367 z"/>
                            </g>
                            <g transform="translate(-1.7, 6.684210526315789)">
                                <path fill="#9be9a8" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#9be9a8" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.3157894736842106 0,1.3157894736842106 z"/>
                                <path fill="#9be9a8" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.3157894736842106 1.7,2.3157894736842106 z"/>
                            </g>
                            <g transform="translate(-3.4, 6.947368421052632)">
                                <path fill="#40c463" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#40c463" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,3.052631578947368 0,2.052631578947368 z"/>
                                <path fill="#40c463" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,2.052631578947368 1.7,3.052631578947368 z"/>
                            </g>
                            <g transform="translate(-5.1, 8.263157894736842)">
                                <path fill="#40c463" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#40c463" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.736842105263158 0,1.736842105263158 z"/>
                                <path fill="#40c463" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.736842105263158 1.7,2.736842105263158 z"/>
                            </g>
                            <g transform="translate(-6.8, 9.578947368421053)">
                                <path fill="#9be9a8" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#9be9a8" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.4210526315789473 0,1.4210526315789473 z"/>
                                <path fill="#9be9a8" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.4210526315789473 1.7,2.4210526315789473 z"/>
                            </g>
                            <g transform="translate(-8.5, 10.368421052631579)">
                                <path fill="#40c463" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#40c463" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.6315789473684212 0,1.631578947368421 z"/>
                                <path fill="#40c463" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.631578947368421 1.7,2.6315789473684212 z"/>
                            </g>
                            <g transform="translate(-10.2, 11.263157894736842)">
                                <path fill="#40c463" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#40c463" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.736842105263158 0,1.736842105263158 z"/>
                                <path fill="#40c463" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.736842105263158 1.7,2.736842105263158 z"/>
                            </g>
                        </g>
                        <g transform="translate(68, 40)">
                            <g transform="translate(0, 5.7894736842105265)">
                                <path fill="#9be9a8" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#9be9a8" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.2105263157894735 0,1.2105263157894737 z"/>
                                <path fill="#9be9a8" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.2105263157894737 1.7,2.2105263157894735 z"/>
                            </g>
                            <g transform="translate(-1.7, 6.578947368421053)">
                                <path fill="#40c463" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#40c463" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.4210526315789473 0,1.4210526315789473 z"/>
                                <path fill="#40c463" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.4210526315789473 1.7,2.4210526315789473 z"/>
                            </g>
                            <g transform="translate(-3.4, 7.473684210526315)">
                                <path fill="#30a14e" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#30a14e" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.526315789473684 0,1.526315789473684 z"/>
                                <path fill="#30a14e" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.526315789473684 1.7,2.526315789473684 z"/>
                            </g>
                            <g transform="translate(-5.1, 8.263157894736842)">
                                <path fill="#216e39" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#216e39" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.736842105263158 0,1.736842105263158 z"/>
                                <path fill="#216e39" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.736842105263158 1.7,2.736842105263158 z"/>
                            </g>
                            <g transform="translate(-6.8, 9.578947368421053)">
                                <path fill="#40c463" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#40c463" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.4210526315789473 0,1.4210526315789473 z"/>
                                <path fill="#40c463" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.4210526315789473 1.7,2.4210526315789473 z"/>
                            </g>
                            <g transform="translate(-8.5, 10.473684210526315)">
                                <path fill="#30a14e" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#30a14e" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.526315789473684 0,1.526315789473684 z"/>
                                <path fill="#30a14e" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.526315789473684 1.7,2.526315789473684 z"/>
                            </g>
                            <g transform="translate(-10.2, 11.894736842105264)">
                                <path fill="#9be9a8" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#9be9a8" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.1052631578947367 0,1.1052631578947367 z"/>
                                <path fill="#9be9a8" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.1052631578947367 1.7,2.1052631578947367 z"/>
                            </g>
                        </g>
                        <g transform="translate(69.7, 41)">
                            <g transform="translate(0, 5.578947368421053)">
                                <path fill="#40c463" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#40c463" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.4210526315789473 0,1.4210526315789473 z"/>
                                <path fill="#40c463" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.4210526315789473 1.7,2.4210526315789473 z"/>
                            </g>
                            <g transform="translate(-1.7, 7)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-3.4, 7.578947368421053)">
                                <path fill="#40c463" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#40c463" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.4210526315789473 0,1.4210526315789473 z"/>
                                <path fill="#40c463" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.4210526315789473 1.7,2.4210526315789473 z"/>
                            </g>
                            <g transform="translate(-5.1, 8.473684210526315)">
                                <path fill="#30a14e" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#30a14e" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.526315789473684 0,1.526315789473684 z"/>
                                <path fill="#30a14e" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.526315789473684 1.7,2.526315789473684 z"/>
                            </g>
                            <g transform="translate(-6.8, 9.68421052631579)">
                                <path fill="#40c463" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#40c463" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.3157894736842106 0,1.3157894736842106 z"/>
                                <path fill="#40c463" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.3157894736842106 1.7,2.3157894736842106 z"/>
                            </g>
                            <g transform="translate(-8.5, 10.789473684210527)">
                                <path fill="#9be9a8" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#9be9a8" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.2105263157894735 0,1.2105263157894737 z"/>
                                <path fill="#9be9a8" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.2105263157894737 1.7,2.2105263157894735 z"/>
                            </g>
                            <g transform="translate(-10.2, 11.473684210526315)">
                                <path fill="#30a14e" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#30a14e" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.526315789473684 0,1.526315789473684 z"/>
                                <path fill="#30a14e" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.526315789473684 1.7,2.526315789473684 z"/>
                            </g>
                        </g>
                        <g transform="translate(71.39999999999999, 42)">
                            <g transform="translate(0, 6)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-1.7, 6.368421052631579)">
                                <path fill="#30a14e" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#30a14e" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.6315789473684212 0,1.631578947368421 z"/>
                                <path fill="#30a14e" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.631578947368421 1.7,2.6315789473684212 z"/>
                            </g>
                            <g transform="translate(-3.4, 7.473684210526315)">
                                <path fill="#30a14e" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#30a14e" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.526315789473684 0,1.526315789473684 z"/>
                                <path fill="#30a14e" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.526315789473684 1.7,2.526315789473684 z"/>
                            </g>
                            <g transform="translate(-5.1, 8.157894736842106)">
                                <path fill="#216e39" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#216e39" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.8421052631578947 0,1.8421052631578947 z"/>
                                <path fill="#216e39" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.8421052631578947 1.7,2.8421052631578947 z"/>
                            </g>
                            <g transform="translate(-6.8, 9.157894736842106)">
                                <path fill="#216e39" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#216e39" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.8421052631578947 0,1.8421052631578947 z"/>
                                <path fill="#216e39" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.8421052631578947 1.7,2.8421052631578947 z"/>
                            </g>
                            <g transform="translate(-8.5, 10.368421052631579)">
                                <path fill="#30a14e" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#30a14e" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.6315789473684212 0,1.631578947368421 z"/>
                                <path fill="#30a14e" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.631578947368421 1.7,2.6315789473684212 z"/>
                            </g>
                            <g transform="translate(-10.2, 11.68421052631579)">
                                <path fill="#40c463" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#40c463" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.3157894736842106 0,1.3157894736842106 z"/>
                                <path fill="#40c463" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.3157894736842106 1.7,2.3157894736842106 z"/>
                            </g>
                        </g>
                        <g transform="translate(73.1, 43)">
                            <g transform="translate(0, 6)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-1.7, 6.473684210526315)">
                                <path fill="#30a14e" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#30a14e" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.526315789473684 0,1.526315789473684 z"/>
                                <path fill="#30a14e" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.526315789473684 1.7,2.526315789473684 z"/>
                            </g>
                            <g transform="translate(-3.4, 7.157894736842105)">
                                <path fill="#216e39" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#216e39" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.8421052631578947 0,1.8421052631578947 z"/>
                                <path fill="#216e39" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.8421052631578947 1.7,2.8421052631578947 z"/>
                            </g>
                            <g transform="translate(-5.1, 8.68421052631579)">
                                <path fill="#40c463" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#40c463" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.3157894736842106 0,1.3157894736842106 z"/>
                                <path fill="#40c463" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.3157894736842106 1.7,2.3157894736842106 z"/>
                            </g>
                            <g transform="translate(-6.8, 9.894736842105264)">
                                <path fill="#9be9a8" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#9be9a8" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.1052631578947367 0,1.1052631578947367 z"/>
                                <path fill="#9be9a8" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.1052631578947367 1.7,2.1052631578947367 z"/>
                            </g>
                            <g transform="translate(-8.5, 10.68421052631579)">
                                <path fill="#40c463" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#40c463" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.3157894736842106 0,1.3157894736842106 z"/>
                                <path fill="#40c463" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.3157894736842106 1.7,2.3157894736842106 z"/>
                            </g>
                            <g transform="translate(-10.2, 12)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                        </g>
                        <g transform="translate(74.8, 44)">
                            <g transform="translate(0, 4.842105263157896)">
                                <path fill="#40c463" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#40c463" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,3.1578947368421053 0,2.1578947368421053 z"/>
                                <path fill="#40c463" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,2.1578947368421053 1.7,3.1578947368421053 z"/>
                            </g>
                            <g transform="translate(-1.7, 6.052631578947368)">
                                <path fill="#40c463" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#40c463" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.9473684210526314 0,1.9473684210526314 z"/>
                                <path fill="#40c463" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.9473684210526314 1.7,2.9473684210526314 z"/>
                            </g>
                            <g transform="translate(-3.4, 6)">
                                <path fill="#30a14e" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#30a14e" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,4 0,3 z"/>
                                <path fill="#30a14e" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,3 1.7,4 z"/>
                            </g>
                            <g transform="translate(-5.1, 8.263157894736842)">
                                <path fill="#40c463" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#40c463" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.736842105263158 0,1.736842105263158 z"/>
                                <path fill="#40c463" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.736842105263158 1.7,2.736842105263158 z"/>
                            </g>
                            <g transform="translate(-6.8, 7.157894736842106)">
                                <path fill="#216e39" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#216e39" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,4.842105263157895 0,3.8421052631578947 z"/>
                                <path fill="#216e39" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,3.8421052631578947 1.7,4.842105263157895 z"/>
                            </g>
                            <g transform="translate(-8.5, 9.947368421052632)">
                                <path fill="#40c463" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#40c463" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,3.052631578947368 0,2.052631578947368 z"/>
                                <path fill="#40c463" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,2.052631578947368 1.7,3.052631578947368 z"/>
                            </g>
                            <g transform="translate(-10.2, 10.736842105263158)">
                                <path fill="#40c463" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#40c463" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,3.263157894736842 0,2.263157894736842 z"/>
                                <path fill="#40c463" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,2.263157894736842 1.7,3.263157894736842 z"/>
                            </g>
                        </g>
                        <g transform="translate(76.5, 45)">
                            <g transform="translate(0, 5.473684210526315)">
                                <path fill="#9be9a8" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#9be9a8" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.526315789473684 0,1.526315789473684 z"/>
                                <path fill="#9be9a8" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.526315789473684 1.7,2.526315789473684 z"/>
                            </g>
                            <g transform="translate(-1.7, 5.947368421052632)">
                                <path fill="#40c463" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#40c463" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,3.052631578947368 0,2.052631578947368 z"/>
                                <path fill="#40c463" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,2.052631578947368 1.7,3.052631578947368 z"/>
                            </g>
                            <g transform="translate(-3.4, 7.7894736842105265)">
                                <path fill="#9be9a8" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#9be9a8" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.2105263157894735 0,1.2105263157894737 z"/>
                                <path fill="#9be9a8" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.2105263157894737 1.7,2.2105263157894735 z"/>
                            </g>
                            <g transform="translate(-5.1, 8.789473684210527)">
                                <path fill="#9be9a8" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#9be9a8" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.2105263157894735 0,1.2105263157894737 z"/>
                                <path fill="#9be9a8" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.2105263157894737 1.7,2.2105263157894735 z"/>
                            </g>
                            <g transform="translate(-6.8, 9.368421052631579)">
                                <path fill="#9be9a8" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#9be9a8" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.6315789473684212 0,1.631578947368421 z"/>
                                <path fill="#9be9a8" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.631578947368421 1.7,2.6315789473684212 z"/>
                            </g>
                            <g transform="translate(-8.5, 10.157894736842106)">
                                <path fill="#40c463" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#40c463" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.8421052631578947 0,1.8421052631578947 z"/>
                                <path fill="#40c463" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.8421052631578947 1.7,2.8421052631578947 z"/>
                            </g>
                            <g transform="translate(-10.2, 11.368421052631579)">
                                <path fill="#9be9a8" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#9be9a8" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.6315789473684212 0,1.631578947368421 z"/>
                                <path fill="#9be9a8" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.631578947368421 1.7,2.6315789473684212 z"/>
                            </g>
                        </g>
                        <g transform="translate(78.2, 46)">
                            <g transform="translate(0, 5.2631578947368425)">
                                <path fill="#40c463" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#40c463" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.736842105263158 0,1.736842105263158 z"/>
                                <path fill="#40c463" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.736842105263158 1.7,2.736842105263158 z"/>
                            </g>
                            <g transform="translate(-1.7, 5.315789473684211)">
                                <path fill="#30a14e" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#30a14e" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,3.6842105263157894 0,2.6842105263157894 z"/>
                                <path fill="#30a14e" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,2.6842105263157894 1.7,3.6842105263157894 z"/>
                            </g>
                            <g transform="translate(-3.4, 6.947368421052632)">
                                <path fill="#40c463" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#40c463" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,3.052631578947368 0,2.052631578947368 z"/>
                                <path fill="#40c463" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,2.052631578947368 1.7,3.052631578947368 z"/>
                            </g>
                            <g transform="translate(-5.1, 8.263157894736842)">
                                <path fill="#40c463" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#40c463" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.736842105263158 0,1.736842105263158 z"/>
                                <path fill="#40c463" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.736842105263158 1.7,2.736842105263158 z"/>
                            </g>
                            <g transform="translate(-6.8, 8.210526315789473)">
                                <path fill="#30a14e" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#30a14e" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,3.789473684210526 0,2.789473684210526 z"/>
                                <path fill="#30a14e" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,2.789473684210526 1.7,3.789473684210526 z"/>
                            </g>
                            <g transform="translate(-8.5, 10.368421052631579)">
                                <path fill="#9be9a8" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#9be9a8" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.6315789473684212 0,1.631578947368421 z"/>
                                <path fill="#9be9a8" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.631578947368421 1.7,2.6315789473684212 z"/>
                            </g>
                            <g transform="translate(-10.2, 11.68421052631579)">
                                <path fill="#9be9a8" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#9be9a8" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.3157894736842106 0,1.3157894736842106 z"/>
                                <path fill="#9be9a8" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.3157894736842106 1.7,2.3157894736842106 z"/>
                            </g>
                        </g>
                        <g transform="translate(79.89999999999999, 47)">
                            <g transform="translate(0, 5.052631578947368)">
                                <path fill="#40c463" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#40c463" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.9473684210526314 0,1.9473684210526314 z"/>
                                <path fill="#40c463" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.9473684210526314 1.7,2.9473684210526314 z"/>
                            </g>
                            <g transform="translate(-1.7, 5.947368421052632)">
                                <path fill="#40c463" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#40c463" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,3.052631578947368 0,2.052631578947368 z"/>
                                <path fill="#40c463" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,2.052631578947368 1.7,3.052631578947368 z"/>
                            </g>
                            <g transform="translate(-3.4, 7.157894736842105)">
                                <path fill="#40c463" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#40c463" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.8421052631578947 0,1.8421052631578947 z"/>
                                <path fill="#40c463" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.8421052631578947 1.7,2.8421052631578947 z"/>
                            </g>
                            <g transform="translate(-5.1, 8.368421052631579)">
                                <path fill="#9be9a8" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#9be9a8" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.6315789473684212 0,1.631578947368421 z"/>
                                <path fill="#9be9a8" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.631578947368421 1.7,2.6315789473684212 z"/>
                            </g>
                            <g transform="translate(-6.8, 10)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-8.5, 10.68421052631579)">
                                <path fill="#9be9a8" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#9be9a8" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.3157894736842106 0,1.3157894736842106 z"/>
                                <path fill="#9be9a8" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.3157894736842106 1.7,2.3157894736842106 z"/>
                            </g>
                            <g transform="translate(-10.2, 11.894736842105264)">
                                <path fill="#9be9a8" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#9be9a8" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.1052631578947367 0,1.1052631578947367 z"/>
                                <path fill="#9be9a8" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.1052631578947367 1.7,2.1052631578947367 z"/>
                            </g>
                        </g>
                        <g transform="translate(81.6, 48)">
                            <g transform="translate(0, 5.684210526315789)">
                                <path fill="#9be9a8" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#9be9a8" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.3157894736842106 0,1.3157894736842106 z"/>
                                <path fill="#9be9a8" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.3157894736842106 1.7,2.3157894736842106 z"/>
                            </g>
                            <g transform="translate(-1.7, 5.631578947368421)">
                                <path fill="#40c463" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#40c463" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,3.3684210526315788 0,2.3684210526315788 z"/>
                                <path fill="#40c463" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,2.3684210526315788 1.7,3.3684210526315788 z"/>
                            </g>
                            <g transform="translate(-3.4, 7.2631578947368425)">
                                <path fill="#9be9a8" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#9be9a8" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.736842105263158 0,1.736842105263158 z"/>
                                <path fill="#9be9a8" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.736842105263158 1.7,2.736842105263158 z"/>
                            </g>
                            <g transform="translate(-5.1, 8.894736842105264)">
                                <path fill="#9be9a8" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#9be9a8" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.1052631578947367 0,1.1052631578947367 z"/>
                                <path fill="#9be9a8" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.1052631578947367 1.7,2.1052631578947367 z"/>
                            </g>
                            <g transform="translate(-6.8, 10)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-8.5, 11)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-10.2, 10.31578947368421)">
                                <path fill="#40c463" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#40c463" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,3.6842105263157894 0,2.6842105263157894 z"/>
                                <path fill="#40c463" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,2.6842105263157894 1.7,3.6842105263157894 z"/>
                            </g>
                        </g>
                        <g transform="translate(83.3, 49)">
                            <g transform="translate(0, 5.052631578947368)">
                                <path fill="#40c463" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#40c463" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.9473684210526314 0,1.9473684210526314 z"/>
                                <path fill="#40c463" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.9473684210526314 1.7,2.9473684210526314 z"/>
                            </g>
                            <g transform="translate(-1.7, 6.2631578947368425)">
                                <path fill="#9be9a8" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#9be9a8" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.736842105263158 0,1.736842105263158 z"/>
                                <path fill="#9be9a8" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.736842105263158 1.7,2.736842105263158 z"/>
                            </g>
                            <g transform="translate(-3.4, 6.842105263157896)">
                                <path fill="#40c463" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#40c463" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,3.1578947368421053 0,2.1578947368421053 z"/>
                                <path fill="#40c463" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,2.1578947368421053 1.7,3.1578947368421053 z"/>
                            </g>
                            <g transform="translate(-5.1, 8.578947368421053)">
                                <path fill="#9be9a8" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#9be9a8" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.4210526315789473 0,1.4210526315789473 z"/>
                                <path fill="#9be9a8" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.4210526315789473 1.7,2.4210526315789473 z"/>
                            </g>
                            <g transform="translate(-6.8, 8.947368421052632)">
                                <path fill="#40c463" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#40c463" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,3.052631578947368 0,2.052631578947368 z"/>
                                <path fill="#40c463" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,2.052631578947368 1.7,3.052631578947368 z"/>
                            </g>
                            <g transform="translate(-8.5, 9.31578947368421)">
                                <path fill="#40c463" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#40c463" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,3.6842105263157894 0,2.6842105263157894 z"/>
                                <path fill="#40c463" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,2.6842105263157894 1.7,3.6842105263157894 z"/>
                            </g>
                            <g transform="translate(-10.2, 11.894736842105264)">
                                <path fill="#9be9a8" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#9be9a8" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.1052631578947367 0,1.1052631578947367 z"/>
                                <path fill="#9be9a8" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.1052631578947367 1.7,2.1052631578947367 z"/>
                            </g>
                        </g>
                        <g transform="translate(85, 50)">
                            <g transform="translate(0, 5.684210526315789)">
                                <path fill="#9be9a8" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#9be9a8" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.3157894736842106 0,1.3157894736842106 z"/>
                                <path fill="#9be9a8" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.3157894736842106 1.7,2.3157894736842106 z"/>
                            </g>
                            <g transform="translate(-1.7, 3.6315789473684212)">
                                <path fill="#216e39" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#216e39" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,5.368421052631579 0,4.368421052631579 z"/>
                                <path fill="#216e39" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,4.368421052631579 1.7,5.368421052631579 z"/>
                            </g>
                            <g transform="translate(-3.4, 6.421052631578948)">
                                <path fill="#40c463" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#40c463" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,3.5789473684210527 0,2.5789473684210527 z"/>
                                <path fill="#40c463" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,2.5789473684210527 1.7,3.5789473684210527 z"/>
                            </g>
                            <g transform="translate(-5.1, 7)">
                                <path fill="#30a14e" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#30a14e" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,4 0,3 z"/>
                                <path fill="#30a14e" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,3 1.7,4 z"/>
                            </g>
                            <g transform="translate(-6.8, 8.842105263157896)">
                                <path fill="#40c463" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#40c463" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,3.1578947368421053 0,2.1578947368421053 z"/>
                                <path fill="#40c463" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,2.1578947368421053 1.7,3.1578947368421053 z"/>
                            </g>
                            <g transform="translate(-8.5, 9.631578947368421)">
                                <path fill="#40c463" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#40c463" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,3.3684210526315788 0,2.3684210526315788 z"/>
                                <path fill="#40c463" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,2.3684210526315788 1.7,3.3684210526315788 z"/>
                            </g>
                            <g transform="translate(-10.2, 11.789473684210527)">
                                <path fill="#9be9a8" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#9be9a8" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.2105263157894735 0,1.2105263157894737 z"/>
                                <path fill="#9be9a8" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.2105263157894737 1.7,2.2105263157894735 z"/>
                            </g>
                        </g>
                        <g transform="translate(86.7, 51)">
                            <g transform="translate(0, 4.842105263157896)">
                                <path fill="#40c463" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#40c463" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,3.1578947368421053 0,2.1578947368421053 z"/>
                                <path fill="#40c463" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,2.1578947368421053 1.7,3.1578947368421053 z"/>
                            </g>
                            <g transform="translate(-1.7, 6.473684210526315)">
                                <path fill="#9be9a8" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#9be9a8" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.526315789473684 0,1.526315789473684 z"/>
                                <path fill="#9be9a8" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.526315789473684 1.7,2.526315789473684 z"/>
                            </g>
                            <g transform="translate(-3.4, 6.315789473684211)">
                                <path fill="#40c463" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#40c463" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,3.6842105263157894 0,2.6842105263157894 z"/>
                                <path fill="#40c463" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,2.6842105263157894 1.7,3.6842105263157894 z"/>
                            </g>
                            <g transform="translate(-5.1, 6.2631578947368425)">
                                <path fill="#216e39" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#216e39" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,4.7368421052631575 0,3.7368421052631575 z"/>
                                <path fill="#216e39" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,3.7368421052631575 1.7,4.7368421052631575 z"/>
                            </g>
                            <g transform="translate(-6.8, 8.526315789473685)">
                                <path fill="#40c463" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#40c463" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,3.473684210526316 0,2.473684210526316 z"/>
                                <path fill="#40c463" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,2.473684210526316 1.7,3.473684210526316 z"/>
                            </g>
                            <g transform="translate(-8.5, 9.631578947368421)">
                                <path fill="#40c463" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#40c463" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,3.3684210526315788 0,2.3684210526315788 z"/>
                                <path fill="#40c463" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,2.3684210526315788 1.7,3.3684210526315788 z"/>
                            </g>
                            <g transform="translate(-10.2, 12)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                        </g>
                        <g transform="translate(88.39999999999999, 52)">
                            <g transform="translate(0, 6)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-1.7, 2.473684210526316)">
                                <path fill="#216e39" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#216e39" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,6.526315789473684 0,5.526315789473684 z"/>
                                <path fill="#216e39" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,5.526315789473684 1.7,6.526315789473684 z"/>
                            </g>
                            <g transform="translate(-3.4, 2)">
                                <path fill="#216e39" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#216e39" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,8 0,7 z"/>
                                <path fill="#216e39" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,7 1.7,8 z"/>
                            </g>
                            <g transform="translate(-5.1, 5.947368421052632)">
                                <path fill="#30a14e" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#30a14e" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,5.052631578947368 0,4.052631578947368 z"/>
                                <path fill="#30a14e" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,4.052631578947368 1.7,5.052631578947368 z"/>
                            </g>
                            <g transform="translate(-6.8, 8.631578947368421)">
                                <path fill="#9be9a8" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#9be9a8" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,3.3684210526315788 0,2.3684210526315788 z"/>
                                <path fill="#9be9a8" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,2.3684210526315788 1.7,3.3684210526315788 z"/>
                            </g>
                            <g transform="translate(-8.5, 9)">
                                <path fill="#40c463" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#40c463" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,4 0,3 z"/>
                                <path fill="#40c463" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,3 1.7,4 z"/>
                            </g>
                            <g transform="translate(-10.2, 11.68421052631579)">
                                <path fill="#9be9a8" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#9be9a8" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.3157894736842106 0,1.3157894736842106 z"/>
                                <path fill="#9be9a8" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.3157894736842106 1.7,2.3157894736842106 z"/>
                            </g>
                        </g>
                    </g>
                </svg>
            </section>
        </div>
        <div xmlns="http://www.w3.org/1999/xhtml" id="metrics-end"></div>
    </foreignObject>
</svg>
